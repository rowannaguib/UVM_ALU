package pkg;
	import uvm_pkg::*;
 	`include "uvm_macros.svh"
	`include "configuration.sv"
	`include "transaction.sv"
	`include "sequence.sv"
	`include "driver.sv"
	`include "monitor_before.sv"
	`include "monitor_after.sv"
	`include "agent.sv"
	`include "scoreboard.sv"
	`include "cov.svh"
	`include "env.sv"
	`include "test.sv"
endpackage: pkg
